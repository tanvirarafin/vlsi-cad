magic
tech sky130A
timestamp 1634854909
<< nwell >>
rect -239 16 50 234
<< nmos >>
rect -91 -113 -75 -71
<< pmos >>
rect -91 63 -76 131
<< ndiff >>
rect -137 -89 -91 -71
rect -137 -106 -126 -89
rect -109 -106 -91 -89
rect -137 -113 -91 -106
rect -75 -88 -39 -71
rect -75 -105 -61 -88
rect -44 -105 -39 -88
rect -75 -113 -39 -105
<< pdiff >>
rect -132 109 -91 131
rect -132 91 -123 109
rect -105 91 -91 109
rect -132 63 -91 91
rect -76 106 -31 131
rect -76 88 -62 106
rect -45 88 -31 106
rect -76 63 -31 88
<< ndiffc >>
rect -126 -106 -109 -89
rect -61 -105 -44 -88
<< pdiffc >>
rect -123 91 -105 109
rect -62 88 -45 106
<< psubdiff >>
rect -189 -157 -147 -145
rect -189 -174 -175 -157
rect -158 -174 -147 -157
rect -189 -187 -147 -174
rect -69 -156 -24 -145
rect -69 -174 -55 -156
rect -37 -174 -24 -156
rect -69 -187 -24 -174
<< nsubdiff >>
rect -179 197 -130 210
rect -179 179 -163 197
rect -145 179 -130 197
rect -63 199 -21 210
rect -63 182 -51 199
rect -34 182 -21 199
rect -179 167 -130 179
rect -63 174 -21 182
<< psubdiffcont >>
rect -175 -174 -158 -157
rect -55 -174 -37 -156
<< nsubdiffcont >>
rect -163 179 -145 197
rect -51 182 -34 199
<< poly >>
rect -91 131 -76 181
rect -91 16 -76 63
rect -91 -11 -75 16
rect -145 -20 -75 -11
rect -145 -38 -135 -20
rect -118 -38 -75 -20
rect -145 -44 -75 -38
rect -91 -71 -75 -44
rect -91 -134 -75 -113
<< polycont >>
rect -135 -38 -118 -20
<< locali >>
rect -180 199 -24 205
rect -180 197 -51 199
rect -180 179 -163 197
rect -145 182 -51 197
rect -34 182 -24 199
rect -145 179 -24 182
rect -180 174 -24 179
rect -131 109 -95 174
rect -131 91 -123 109
rect -105 91 -95 109
rect -131 84 -95 91
rect -69 106 -34 121
rect -69 88 -62 106
rect -45 88 -34 106
rect -131 81 -96 84
rect -179 -20 -109 -11
rect -179 -38 -135 -20
rect -118 -38 -109 -20
rect -179 -45 -109 -38
rect -135 -89 -100 -79
rect -135 -106 -126 -89
rect -109 -106 -100 -89
rect -135 -145 -100 -106
rect -69 -88 -34 88
rect -69 -105 -61 -88
rect -44 -105 -34 -88
rect -69 -112 -34 -105
rect -190 -156 -20 -145
rect -190 -157 -55 -156
rect -190 -174 -175 -157
rect -158 -174 -55 -157
rect -37 -174 -20 -156
rect -190 -187 -20 -174
rect -188 -192 -20 -187
<< labels >>
rlabel locali -163 -27 -163 -27 1 in
rlabel locali -46 -24 -46 -24 1 out
rlabel locali -91 198 -91 198 1 vdd
rlabel locali -118 -167 -118 -167 1 gnd
<< end >>
