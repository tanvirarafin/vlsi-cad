* NGSPICE file created from inverter.ext - technology: sky130A


* Top level circuit inverter

X0 out in gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=160000u
X1 out in vdd vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=680000u l=150000u
C0 out in 0.03fF
C1 out vdd 0.08fF
C2 vdd in 0.03fF
C3 out gnd 0.21fF
C4 in gnd 0.44fF
C5 vdd gnd 0.89fF
.end

