`timescale 1ns/1ns
module example_4_simple_mips;
endmodule
	
